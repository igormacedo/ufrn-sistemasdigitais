library verilog;
use verilog.vl_types.all;
entity TestLatch_vlg_check_tst is
    port(
        \OUt\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TestLatch_vlg_check_tst;
