-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: altfp_convert1.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" OPERATION="INT2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=19 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=19 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:33:SJ cbx_altfp_convert 2013:06:12:18:03:33:SJ cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_altsyncram 2013:06:12:18:03:33:SJ cbx_cycloneii 2013:06:12:18:03:33:SJ cbx_lpm_abs 2013:06:12:18:03:33:SJ cbx_lpm_add_sub 2013:06:12:18:03:33:SJ cbx_lpm_compare 2013:06:12:18:03:33:SJ cbx_lpm_decode 2013:06:12:18:03:33:SJ cbx_lpm_divide 2013:06:12:18:03:33:SJ cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ cbx_stratix 2013:06:12:18:03:33:SJ cbx_stratixii 2013:06:12:18:03:33:SJ cbx_stratixiii 2013:06:12:18:03:33:SJ cbx_stratixv 2013:06:12:18:03:33:SJ cbx_util_mgl 2013:06:12:18:03:33:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone II" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=19 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 13.0 cbx_altbarrel_shift 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = reg 42 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altbarrel_shift_grf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (18 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (18 DOWNTO 0)
	 ); 
 END altfp_convert1_altbarrel_shift_grf;

 ARCHITECTURE RTL OF altfp_convert1_altbarrel_shift_grf IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(18 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(18 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w53w54w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w74w75w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w123w124w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w118w119w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w142w143w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w137w138w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w48w49w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w69w70w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w113w114w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w132w133w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range112w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range112w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range131w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range131w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range110w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range129w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range46w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range67w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range112w113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range112w123w124w125w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range131w142w143w144w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w104w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w126w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w145w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (113 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (94 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w117w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w121w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w136w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w140w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range50w_w_w_sbit_w_range41w_range51w52w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range71w_w_w_sbit_w_range64w_range72w73w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range55w_w_pad_w_range50w56w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range76w_w_pad_w_range71w77w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range41w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range64w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range84w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range106w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range128w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range105w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range146w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range55w_w_pad_w_range50w56w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w53w54w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w53w(0) AND wire_altbarrel_shift5_w_w_pad_w_range50w_w_w_sbit_w_range41w_range51w52w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range76w_w_pad_w_range71w77w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w74w75w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w74w(0) AND wire_altbarrel_shift5_w_w_pad_w_range71w_w_w_sbit_w_range64w_range72w73w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w(0) AND wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w123w124w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range112w123w(0) AND wire_altbarrel_shift5_w121w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w118w119w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range112w118w(0) AND wire_altbarrel_shift5_w117w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w142w143w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range131w142w(0) AND wire_altbarrel_shift5_w140w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w137w138w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range131w137w(0) AND wire_altbarrel_shift5_w136w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w48w49w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range46w48w(0) AND wire_altbarrel_shift5_w_sbit_w_range41w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w69w70w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range67w69w(0) AND wire_altbarrel_shift5_w_sbit_w_range64w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w(0) AND wire_altbarrel_shift5_w_sbit_w_range84w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w113w114w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range112w113w(0) AND wire_altbarrel_shift5_w_sbit_w_range106w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w132w133w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range131w132w(0) AND wire_altbarrel_shift5_w_sbit_w_range128w(i);
	END GENERATE loop14;
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w58w(0) <= wire_altbarrel_shift5_w_sel_w_range46w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w53w(0) <= wire_altbarrel_shift5_w_sel_w_range46w(0) AND wire_altbarrel_shift5_w_dir_w_range43w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w79w(0) <= wire_altbarrel_shift5_w_sel_w_range67w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w74w(0) <= wire_altbarrel_shift5_w_sel_w_range67w(0) AND wire_altbarrel_shift5_w_dir_w_range65w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w101w(0) <= wire_altbarrel_shift5_w_sel_w_range89w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w96w(0) <= wire_altbarrel_shift5_w_sel_w_range89w(0) AND wire_altbarrel_shift5_w_dir_w_range86w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range112w123w(0) <= wire_altbarrel_shift5_w_sel_w_range112w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range110w122w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range112w118w(0) <= wire_altbarrel_shift5_w_sel_w_range112w(0) AND wire_altbarrel_shift5_w_dir_w_range110w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range131w142w(0) <= wire_altbarrel_shift5_w_sel_w_range131w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range129w141w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range131w137w(0) <= wire_altbarrel_shift5_w_sel_w_range131w(0) AND wire_altbarrel_shift5_w_dir_w_range129w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range43w57w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range43w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range65w78w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range65w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range86w100w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range86w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range110w122w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range110w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range129w141w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range129w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range46w48w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range46w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range67w69w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range67w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range89w91w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range89w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range112w113w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range112w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range131w132w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range131w(0);
	loop15 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w58w59w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w53w54w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w79w80w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w74w75w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w101w102w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w96w97w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range112w123w124w125w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w123w124w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w118w119w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range131w142w143w144w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w142w143w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w137w138w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range46w48w49w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range67w69w70w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w104w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range89w101w102w103w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range89w91w92w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w126w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range112w123w124w125w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range112w113w114w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 18 GENERATE 
		wire_altbarrel_shift5_w145w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range131w142w143w144w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range131w132w133w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(1) & dir_w(3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(113 DOWNTO 95);
	sbit_w <= ( sbit_piper2d & smux_w(75 DOWNTO 57) & sbit_piper1d & smux_w(37 DOWNTO 0) & data);
	sel_w <= ( sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift5_w145w & wire_altbarrel_shift5_w126w & wire_altbarrel_shift5_w104w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range67w79w80w81w82w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range46w58w59w60w61w);
	wire_altbarrel_shift5_w117w <= ( pad_w(7 DOWNTO 0) & sbit_w(75 DOWNTO 65));
	wire_altbarrel_shift5_w121w <= ( sbit_w(67 DOWNTO 57) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift5_w136w <= ( pad_w(15 DOWNTO 0) & sbit_w(94 DOWNTO 92));
	wire_altbarrel_shift5_w140w <= ( sbit_w(78 DOWNTO 76) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift5_w_w_pad_w_range50w_w_w_sbit_w_range41w_range51w52w <= ( pad_w(0) & sbit_w(18 DOWNTO 1));
	wire_altbarrel_shift5_w_w_pad_w_range71w_w_w_sbit_w_range64w_range72w73w <= ( pad_w(1 DOWNTO 0) & sbit_w(37 DOWNTO 21));
	wire_altbarrel_shift5_w_w_pad_w_range93w_w_w_sbit_w_range84w_range94w95w <= ( pad_w(3 DOWNTO 0) & sbit_w(56 DOWNTO 42));
	wire_altbarrel_shift5_w_w_w_sbit_w_range41w_range55w_w_pad_w_range50w56w <= ( sbit_w(17 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift5_w_w_w_sbit_w_range64w_range76w_w_pad_w_range71w77w <= ( sbit_w(35 DOWNTO 19) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift5_w_w_w_sbit_w_range84w_range98w_w_pad_w_range93w99w <= ( sbit_w(52 DOWNTO 38) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift5_w_dir_w_range43w(0) <= dir_w(0);
	wire_altbarrel_shift5_w_dir_w_range65w(0) <= dir_w(1);
	wire_altbarrel_shift5_w_dir_w_range86w(0) <= dir_w(2);
	wire_altbarrel_shift5_w_dir_w_range110w(0) <= dir_w(3);
	wire_altbarrel_shift5_w_dir_w_range129w(0) <= dir_w(4);
	wire_altbarrel_shift5_w_sbit_w_range41w <= sbit_w(18 DOWNTO 0);
	wire_altbarrel_shift5_w_sbit_w_range64w <= sbit_w(37 DOWNTO 19);
	wire_altbarrel_shift5_w_sbit_w_range84w <= sbit_w(56 DOWNTO 38);
	wire_altbarrel_shift5_w_sbit_w_range106w <= sbit_w(75 DOWNTO 57);
	wire_altbarrel_shift5_w_sbit_w_range128w <= sbit_w(94 DOWNTO 76);
	wire_altbarrel_shift5_w_sel_w_range46w(0) <= sel_w(0);
	wire_altbarrel_shift5_w_sel_w_range67w(0) <= sel_w(1);
	wire_altbarrel_shift5_w_sel_w_range89w(0) <= sel_w(2);
	wire_altbarrel_shift5_w_sel_w_range112w(0) <= sel_w(3);
	wire_altbarrel_shift5_w_sel_w_range131w(0) <= sel_w(4);
	wire_altbarrel_shift5_w_smux_w_range105w <= smux_w(56 DOWNTO 38);
	wire_altbarrel_shift5_w_smux_w_range146w <= smux_w(94 DOWNTO 76);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(4) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift5_w_smux_w_range105w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift5_w_smux_w_range146w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --altfp_convert1_altbarrel_shift_grf


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END altfp_convert1_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --altfp_convert1_altpriority_encoder_3v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert1_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --altfp_convert1_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END altfp_convert1_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert1_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder13_w_lg_zero180w & wire_altpriority_encoder13_w_lg_w_lg_zero182w183w);
	altpriority_encoder12 :  altfp_convert1_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder12_q
	  );
	wire_altpriority_encoder13_w_lg_w_lg_zero180w181w(0) <= wire_altpriority_encoder13_w_lg_zero180w(0) AND wire_altpriority_encoder13_q(0);
	wire_altpriority_encoder13_w_lg_zero182w(0) <= wire_altpriority_encoder13_zero AND wire_altpriority_encoder12_q(0);
	wire_altpriority_encoder13_w_lg_zero180w(0) <= NOT wire_altpriority_encoder13_zero;
	wire_altpriority_encoder13_w_lg_w_lg_zero182w183w(0) <= wire_altpriority_encoder13_w_lg_zero182w(0) OR wire_altpriority_encoder13_w_lg_w_lg_zero180w181w(0);
	altpriority_encoder13 :  altfp_convert1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert1_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero198w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero200w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder15_w_lg_zero198w & wire_altpriority_encoder15_w_lg_w_lg_zero200w201w);
	zero <= (wire_altpriority_encoder14_zero AND wire_altpriority_encoder15_zero);
	altpriority_encoder14 :  altfp_convert1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );
	wire_altpriority_encoder15_w_lg_w_lg_zero198w199w(0) <= wire_altpriority_encoder15_w_lg_zero198w(0) AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder15_w_lg_zero200w(0) <= wire_altpriority_encoder15_zero AND wire_altpriority_encoder14_q(0);
	wire_altpriority_encoder15_w_lg_zero198w(0) <= NOT wire_altpriority_encoder15_zero;
	wire_altpriority_encoder15_w_lg_w_lg_zero200w201w(0) <= wire_altpriority_encoder15_w_lg_zero200w(0) OR wire_altpriority_encoder15_w_lg_w_lg_zero198w199w(0);
	altpriority_encoder15 :  altfp_convert1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END altfp_convert1_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero171w172w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero173w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero173w174w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert1_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder11_w_lg_zero171w & wire_altpriority_encoder11_w_lg_w_lg_zero173w174w);
	altpriority_encoder10 :  altfp_convert1_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder10_q
	  );
	loop25 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero171w172w(i) <= wire_altpriority_encoder11_w_lg_zero171w(0) AND wire_altpriority_encoder11_q(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder11_w_lg_zero173w(i) <= wire_altpriority_encoder11_zero AND wire_altpriority_encoder10_q(i);
	END GENERATE loop26;
	wire_altpriority_encoder11_w_lg_zero171w(0) <= NOT wire_altpriority_encoder11_zero;
	loop27 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero173w174w(i) <= wire_altpriority_encoder11_w_lg_zero173w(i) OR wire_altpriority_encoder11_w_lg_w_lg_zero171w172w(i);
	END GENERATE loop27;
	altpriority_encoder11 :  altfp_convert1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert1_altpriority_encoder_be8;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero208w209w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero210w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero210w211w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder17_w_lg_zero208w & wire_altpriority_encoder17_w_lg_w_lg_zero210w211w);
	zero <= (wire_altpriority_encoder16_zero AND wire_altpriority_encoder17_zero);
	altpriority_encoder16 :  altfp_convert1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );
	loop28 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder17_w_lg_w_lg_zero208w209w(i) <= wire_altpriority_encoder17_w_lg_zero208w(0) AND wire_altpriority_encoder17_q(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder17_w_lg_zero210w(i) <= wire_altpriority_encoder17_zero AND wire_altpriority_encoder16_q(i);
	END GENERATE loop29;
	wire_altpriority_encoder17_w_lg_zero208w(0) <= NOT wire_altpriority_encoder17_zero;
	loop30 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder17_w_lg_w_lg_zero210w211w(i) <= wire_altpriority_encoder17_w_lg_zero210w(i) OR wire_altpriority_encoder17_w_lg_w_lg_zero208w209w(i);
	END GENERATE loop30;
	altpriority_encoder17 :  altfp_convert1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder17_q,
		zero => wire_altpriority_encoder17_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END altfp_convert1_altpriority_encoder_r08;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero162w163w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero164w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero164w165w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert1_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder9_w_lg_zero162w & wire_altpriority_encoder9_w_lg_w_lg_zero164w165w);
	altpriority_encoder8 :  altfp_convert1_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder8_q
	  );
	loop31 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero162w163w(i) <= wire_altpriority_encoder9_w_lg_zero162w(0) AND wire_altpriority_encoder9_q(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder9_w_lg_zero164w(i) <= wire_altpriority_encoder9_zero AND wire_altpriority_encoder8_q(i);
	END GENERATE loop32;
	wire_altpriority_encoder9_w_lg_zero162w(0) <= NOT wire_altpriority_encoder9_zero;
	loop33 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero164w165w(i) <= wire_altpriority_encoder9_w_lg_zero164w(i) OR wire_altpriority_encoder9_w_lg_w_lg_zero162w163w(i);
	END GENERATE loop33;
	altpriority_encoder9 :  altfp_convert1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder9_q,
		zero => wire_altpriority_encoder9_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 13.0 cbx_altpriority_encoder 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END altfp_convert1_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero218w219w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero220w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero220w221w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder19_w_lg_zero218w & wire_altpriority_encoder19_w_lg_w_lg_zero220w221w);
	zero <= (wire_altpriority_encoder18_zero AND wire_altpriority_encoder19_zero);
	altpriority_encoder18 :  altfp_convert1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero218w219w(i) <= wire_altpriority_encoder19_w_lg_zero218w(0) AND wire_altpriority_encoder19_q(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder19_w_lg_zero220w(i) <= wire_altpriority_encoder19_zero AND wire_altpriority_encoder18_q(i);
	END GENERATE loop35;
	wire_altpriority_encoder19_w_lg_zero218w(0) <= NOT wire_altpriority_encoder19_zero;
	loop36 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero220w221w(i) <= wire_altpriority_encoder19_w_lg_zero220w(i) OR wire_altpriority_encoder19_w_lg_w_lg_zero218w219w(i);
	END GENERATE loop36;
	altpriority_encoder19 :  altfp_convert1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder19_q,
		zero => wire_altpriority_encoder19_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END altfp_convert1_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF altfp_convert1_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero153w154w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero155w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero155w156w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_zero	:	STD_LOGIC;
	 COMPONENT  altfp_convert1_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert1_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder7_w_lg_zero153w & wire_altpriority_encoder7_w_lg_w_lg_zero155w156w);
	altpriority_encoder6 :  altfp_convert1_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder6_q
	  );
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero153w154w(i) <= wire_altpriority_encoder7_w_lg_zero153w(0) AND wire_altpriority_encoder7_q(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder7_w_lg_zero155w(i) <= wire_altpriority_encoder7_zero AND wire_altpriority_encoder6_q(i);
	END GENERATE loop38;
	wire_altpriority_encoder7_w_lg_zero153w(0) <= NOT wire_altpriority_encoder7_zero;
	loop39 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero155w156w(i) <= wire_altpriority_encoder7_w_lg_zero155w(i) OR wire_altpriority_encoder7_w_lg_w_lg_zero153w154w(i);
	END GENERATE loop39;
	altpriority_encoder7 :  altfp_convert1_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder7_q,
		zero => wire_altpriority_encoder7_zero
	  );

 END RTL; --altfp_convert1_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 2 lpm_compare 1 reg 168 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altfp_convert1_altfp_convert_dtm IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (18 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END altfp_convert1_altfp_convert_dtm;

 ARCHITECTURE RTL OF altfp_convert1_altfp_convert_dtm IS

	 SIGNAL  wire_altbarrel_shift5_data	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(17 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(17 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_w_lg_alb22w23w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb21w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cmpr4_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector18w19w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  priority_pad_one_w :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 COMPONENT  altfp_convert1_altbarrel_shift_grf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(18 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(18 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altfp_convert1_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop40 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector18w19w(i) <= wire_w_lg_max_neg_value_selector18w(0) AND exponent_zero_w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 17 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_max_neg_value_selector17w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 17 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop43;
	wire_w_lg_max_neg_value_selector18w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	aclr <= '0';
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10010000";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector18w19w OR wire_w_lg_max_neg_value_selector17w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_cmpr4_w_lg_w_lg_alb22w23w OR wire_cmpr4_w_lg_alb21w);
	exponent_output_w <= wire_add_sub3_result;
	exponent_rounded <= exponent_bus_pre_reg;
	exponent_zero_w <= (OTHERS => '0');
	int_a <= dataa(17 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(22 DOWNTO 0);
	mantissa_pre_round <= ( shifted_mag_int_a(17 DOWNTO 0) & "000000");
	mantissa_rounded <= mantissa_pre_round_reg;
	max_neg_value_selector <= (wire_cmpr4_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10010001";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	priority_pad_one_w <= (OTHERS => '1');
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	shifted_mag_int_a <= wire_altbarrel_shift5_result(17 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(18);
	zero_padding_w <= (OTHERS => '0');
	wire_altbarrel_shift5_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift5 :  altfp_convert1_altbarrel_shift_grf
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift5_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift5_result
	  );
	wire_altpriority_encoder2_data <= ( prio_mag_int_a & priority_pad_one_w);
	altpriority_encoder2 :  altfp_convert1_altpriority_encoder_qb6
	  PORT MAP ( 
		data => wire_altpriority_encoder2_data,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "000000000000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 18,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_add_sub3_result
	  );
	loop44 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_w_lg_alb22w23w(i) <= wire_cmpr4_w_lg_alb22w(0) AND exponent_output_w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_alb21w(i) <= wire_cmpr4_alb AND exceptions_value(i);
	END GENERATE loop45;
	wire_cmpr4_w_lg_alb22w(0) <= NOT wire_cmpr4_alb;
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr4_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --altfp_convert1_altfp_convert_dtm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altfp_convert1 IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (18 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END altfp_convert1;


ARCHITECTURE RTL OF altfp_convert1 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT altfp_convert1_altfp_convert_dtm
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (18 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	altfp_convert1_altfp_convert_dtm_component : altfp_convert1_altfp_convert_dtm
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "INT2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "19"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "19"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 19 0 INPUT NODEFVAL "dataa[18..0]"
-- Retrieval info: CONNECT: @dataa 0 0 19 0 dataa 0 0 19 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altfp_convert1.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
