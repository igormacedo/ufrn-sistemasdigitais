library verilog;
use verilog.vl_types.all;
entity rising_edge_detector_vlg_vec_tst is
end rising_edge_detector_vlg_vec_tst;
