library verilog;
use verilog.vl_types.all;
entity controller_block_vlg_vec_tst is
end controller_block_vlg_vec_tst;
