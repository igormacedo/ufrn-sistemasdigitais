library verilog;
use verilog.vl_types.all;
entity controlecooler_vlg_vec_tst is
end controlecooler_vlg_vec_tst;
