library verilog;
use verilog.vl_types.all;
entity TestLatch_vlg_vec_tst is
end TestLatch_vlg_vec_tst;
