library verilog;
use verilog.vl_types.all;
entity dflipflop_vlg_vec_tst is
end dflipflop_vlg_vec_tst;
